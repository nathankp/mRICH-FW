------------------------------------------------------------------------------
--   ____  ____
--  /   /\/   /
-- /___/  \  /    Vendor: Xilinx
-- \   \   \/     Version : 1.11
--  \   \         Application : Spartan-6 FPGA GTP Transceiver Wizard
--  /   /         Filename : pcs_pma_s6_gtpwizard_top.vhd
-- /___/   /\       
-- \   \  /  \ 
--  \___\/\___\
--
--
-- Module PCS_PMA_S6_GTPWIZARD_TOP
-- Generated by Xilinx Spartan-6 FPGA GTP Transceiver Wizard
-- 
-- 
-- (c) Copyright 2009 - 2011 Xilinx, Inc. All rights reserved.
-- 
-- This file contains confidential and proprietary information
-- of Xilinx, Inc. and is protected under U.S. and
-- international copyright and other intellectual property
-- laws.
-- 
-- DISCLAIMER
-- This disclaimer is not a license and does not grant any
-- rights to the materials distributed herewith. Except as
-- otherwise provided in a valid license issued to you by
-- Xilinx, and to the maximum extent permitted by applicable
-- law: (1) THESE MATERIALS ARE MADE AVAILABLE "AS IS" AND
-- WITH ALL FAULTS, AND XILINX HEREBY DISCLAIMS ALL WARRANTIES
-- AND CONDITIONS, EXPRESS, IMPLIED, OR STATUTORY, INCLUDING
-- BUT NOT LIMITED TO WARRANTIES OF MERCHANTABILITY, NON-
-- INFRINGEMENT, OR FITNESS FOR ANY PARTICULAR PURPOSE; and
-- (2) Xilinx shall not be liable (whether in contract or tort,
-- including negligence, or under any other theory of
-- liability) for any loss or damage of any kind or nature
-- related to, arising under or in connection with these
-- materials, including for any direct, or any indirect,
-- special, incidental, or consequential loss or damage
-- (including loss of data, profits, goodwill, or any type of
-- loss or damage suffered as a result of any action brought
-- by a third party) even if such damage or loss was
-- reasonably foreseeable or Xilinx had been advised of the
-- possibility of the same.
-- 
-- CRITICAL APPLICATIONS
-- Xilinx products are not designed or intended to be fail-
-- safe, or for use in any application requiring fail-safe
-- performance, such as life-support or safety devices or
-- systems, Class III medical devices, nuclear facilities,
-- applications related to the deployment of airbags, or any
-- other applications that could lead to death, personal
-- injury, or severe property or environmental damage
-- (individually and collectively, "Critical
-- Applications"). Customer assumes the sole risk and
-- liability of any use of Xilinx products in Critical
-- Applications, subject only to applicable laws and
-- regulations governing limitations on product liability.
-- 
-- THIS COPYRIGHT NOTICE AND DISCLAIMER MUST BE RETAINED AS
-- PART OF THIS FILE AT ALL TIMES. 


library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library UNISIM;
use UNISIM.VCOMPONENTS.ALL;



--***********************************Entity Declaration************************

entity pcs_pma_s6_gtpwizard_top is
generic
(
    EXAMPLE_CONFIG_INDEPENDENT_LANES        : integer   := 1;
    EXAMPLE_LANE_WITH_START_CHAR            : integer   := 0;
    EXAMPLE_WORDS_IN_BRAM                   : integer   := 512;
    EXAMPLE_SIM_GTPRESET_SPEEDUP            : integer   := 0;
    EXAMPLE_USE_CHIPSCOPE                   : integer   := 1;     -- Set to 1 to use Chipscope to drive resets
    EXAMPLE_SIMULATION                      : integer   := 0     -- Set to 1 in testbench for simulation
);
port
(
    TILE0_GTP0_REFCLK_PAD_N_IN              : in   std_logic;
    TILE0_GTP0_REFCLK_PAD_P_IN              : in   std_logic;
    GTP0_RESET_IN                           : in   std_logic;
    GTP1_RESET_IN                           : in   std_logic;
    TILE0_GTP0_PLLLKDET_OUT                 : out  std_logic;
    TRACK_DATA_OUT                          : out  std_logic;
    RXN_IN                                  : in   std_logic_vector(1 downto 0);
    RXP_IN                                  : in   std_logic_vector(1 downto 0);
    TXN_OUT                                 : out  std_logic_vector(1 downto 0);
    TXP_OUT                                 : out  std_logic_vector(1 downto 0)
);
end pcs_pma_s6_gtpwizard_top;
    
architecture RTL of pcs_pma_s6_gtpwizard_top is

--**************************Component Declarations*****************************


component pcs_pma_s6_gtpwizard 
generic
(
    -- Simulation attributes  
    WRAPPER_SIM_GTPRESET_SPEEDUP    : integer   := 0; -- Set to 1 to speed up sim reset
    WRAPPER_CLK25_DIVIDER_0         : integer   := 4;
    WRAPPER_CLK25_DIVIDER_1         : integer   := 4;
    WRAPPER_PLL_DIVSEL_FB_0         : integer   := 5;
    WRAPPER_PLL_DIVSEL_FB_1         : integer   := 5;
    WRAPPER_PLL_DIVSEL_REF_0        : integer   := 2;
    WRAPPER_PLL_DIVSEL_REF_1        : integer   := 2;
    WRAPPER_SIMULATION              : integer   := 0  -- Set to 1 for simulation  
);
port
(
    
    --_________________________________________________________________________
    --_________________________________________________________________________
    --TILE0  (X0_Y0)

 
    ------------------------ Loopback and Powerdown Ports ----------------------
    TILE0_LOOPBACK0_IN                      : in   std_logic_vector(2 downto 0);
    TILE0_LOOPBACK1_IN                      : in   std_logic_vector(2 downto 0);
    TILE0_RXPOWERDOWN0_IN                   : in   std_logic_vector(1 downto 0);
    TILE0_RXPOWERDOWN1_IN                   : in   std_logic_vector(1 downto 0);
    TILE0_TXPOWERDOWN0_IN                   : in   std_logic_vector(1 downto 0);
    TILE0_TXPOWERDOWN1_IN                   : in   std_logic_vector(1 downto 0);
    --------------------------------- PLL Ports --------------------------------
    TILE0_CLK00_IN                          : in   std_logic;
    TILE0_CLK01_IN                          : in   std_logic;
    TILE0_GTPRESET0_IN                      : in   std_logic;
    TILE0_GTPRESET1_IN                      : in   std_logic;
    TILE0_PLLLKDET0_OUT                     : out  std_logic;
    TILE0_RESETDONE0_OUT                    : out  std_logic;
    TILE0_RESETDONE1_OUT                    : out  std_logic;
    ----------------------- Receive Ports - 8b10b Decoder ----------------------
    TILE0_RXCHARISCOMMA0_OUT                : out  std_logic;
    TILE0_RXCHARISCOMMA1_OUT                : out  std_logic;
    TILE0_RXCHARISK0_OUT                    : out  std_logic;
    TILE0_RXCHARISK1_OUT                    : out  std_logic;
    TILE0_RXDISPERR0_OUT                    : out  std_logic;
    TILE0_RXDISPERR1_OUT                    : out  std_logic;
    TILE0_RXNOTINTABLE0_OUT                 : out  std_logic;
    TILE0_RXNOTINTABLE1_OUT                 : out  std_logic;
    TILE0_RXRUNDISP0_OUT                    : out  std_logic;
    TILE0_RXRUNDISP1_OUT                    : out  std_logic;
    ---------------------- Receive Ports - Clock Correction --------------------
    TILE0_RXCLKCORCNT0_OUT                  : out  std_logic_vector(2 downto 0);
    TILE0_RXCLKCORCNT1_OUT                  : out  std_logic_vector(2 downto 0);
    --------------- Receive Ports - Comma Detection and Alignment --------------
    TILE0_RXENMCOMMAALIGN0_IN               : in   std_logic;
    TILE0_RXENMCOMMAALIGN1_IN               : in   std_logic;
    TILE0_RXENPCOMMAALIGN0_IN               : in   std_logic;
    TILE0_RXENPCOMMAALIGN1_IN               : in   std_logic;
    ------------------- Receive Ports - RX Data Path interface -----------------
    TILE0_RXDATA0_OUT                       : out  std_logic_vector(7 downto 0);
    TILE0_RXDATA1_OUT                       : out  std_logic_vector(7 downto 0);
    TILE0_RXRECCLK0_OUT                     : out  std_logic;
    TILE0_RXRECCLK1_OUT                     : out  std_logic;
    TILE0_RXRESET0_IN                       : in   std_logic;
    TILE0_RXRESET1_IN                       : in   std_logic;
    TILE0_RXUSRCLK0_IN                      : in   std_logic;
    TILE0_RXUSRCLK1_IN                      : in   std_logic;
    TILE0_RXUSRCLK20_IN                     : in   std_logic;
    TILE0_RXUSRCLK21_IN                     : in   std_logic;
    ------- Receive Ports - RX Driver,OOB signalling,Coupling and Eq.,CDR ------
    TILE0_RXN0_IN                           : in   std_logic;
    TILE0_RXN1_IN                           : in   std_logic;
    TILE0_RXP0_IN                           : in   std_logic;
    TILE0_RXP1_IN                           : in   std_logic;
    ----------- Receive Ports - RX Elastic Buffer and Phase Alignment ----------
    TILE0_RXBUFRESET0_IN                    : in   std_logic;
    TILE0_RXBUFRESET1_IN                    : in   std_logic;
    TILE0_RXBUFSTATUS0_OUT                  : out  std_logic_vector(2 downto 0);
    TILE0_RXBUFSTATUS1_OUT                  : out  std_logic_vector(2 downto 0);
    ---------------------------- TX/RX Datapath Ports --------------------------
    TILE0_GTPCLKOUT0_OUT                    : out  std_logic_vector(1 downto 0);
    TILE0_GTPCLKOUT1_OUT                    : out  std_logic_vector(1 downto 0);
    ------------------- Transmit Ports - 8b10b Encoder Control -----------------
    TILE0_TXCHARDISPMODE0_IN                : in   std_logic;
    TILE0_TXCHARDISPMODE1_IN                : in   std_logic;
    TILE0_TXCHARDISPVAL0_IN                 : in   std_logic;
    TILE0_TXCHARDISPVAL1_IN                 : in   std_logic;
    TILE0_TXCHARISK0_IN                     : in   std_logic;
    TILE0_TXCHARISK1_IN                     : in   std_logic;
    --------------- Transmit Ports - TX Buffer and Phase Alignment -------------
    TILE0_TXBUFSTATUS0_OUT                  : out  std_logic_vector(1 downto 0);
    TILE0_TXBUFSTATUS1_OUT                  : out  std_logic_vector(1 downto 0);
    ------------------ Transmit Ports - TX Data Path interface -----------------
    TILE0_TXDATA0_IN                        : in   std_logic_vector(7 downto 0);
    TILE0_TXDATA1_IN                        : in   std_logic_vector(7 downto 0);
    TILE0_TXOUTCLK0_OUT                     : out  std_logic;
    TILE0_TXOUTCLK1_OUT                     : out  std_logic;
    TILE0_TXRESET0_IN                       : in   std_logic;
    TILE0_TXRESET1_IN                       : in   std_logic;
    TILE0_TXUSRCLK0_IN                      : in   std_logic;
    TILE0_TXUSRCLK1_IN                      : in   std_logic;
    TILE0_TXUSRCLK20_IN                     : in   std_logic;
    TILE0_TXUSRCLK21_IN                     : in   std_logic;
    --------------- Transmit Ports - TX Driver and OOB signalling --------------
    TILE0_TXN0_OUT                          : out  std_logic;
    TILE0_TXN1_OUT                          : out  std_logic;
    TILE0_TXP0_OUT                          : out  std_logic;
    TILE0_TXP1_OUT                          : out  std_logic


);
end component;


component MGT_USRCLK_SOURCE 
generic
(
    FREQUENCY_MODE   : string   := "LOW";
    DIVIDE_2         : boolean  := false;    
    FEEDBACK         : string   := "1X";
    DIVIDE           : real     := 2.0    
);
port
(
    DIV1_OUT                : out std_logic;
    DIV2_OUT                : out std_logic;
    CLK2X_OUT               : out std_logic;
    DCM_LOCKED_OUT          : out std_logic;
    CLK_IN                  : in  std_logic;
    FB_IN                   : in  std_logic;
    DCM_RESET_IN            : in  std_logic

);
end component;

component FRAME_GEN 
generic
(
    WORDS_IN_BRAM : integer    :=   256;
    MEM_00       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_01       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_02       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_03       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_04       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_05       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_06       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_07       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_08       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_09       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_0A       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_0B       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_0C       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_0D       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_0E       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_0F       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_10       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_11       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_12       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_13       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_14       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_15       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_16       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_17       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_18       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_19       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_1A       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_1B       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_1C       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_1D       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_1E       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_1F       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_20       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_21       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_22       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_23       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_24       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_25       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_26       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_27       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_28       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_29       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_2A       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_2B       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_2C       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_2D       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_2E       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_2F       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_30       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_31       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_32       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_33       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_34       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_35       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_36       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_37       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_38       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_39       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_3A       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_3B       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_3C       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_3D       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_3E       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_3F       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEMP_00      : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEMP_01      : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEMP_02      : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEMP_03      : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEMP_04      : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEMP_05      : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEMP_06      : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEMP_07      : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000"
);    
port
(
    -- User Interface
    TX_DATA             : out   std_logic_vector(39 downto 0);
    TX_CHARISK          : out   std_logic_vector(3 downto 0); 

    -- System Interface
    USER_CLK            : in    std_logic;
    SYSTEM_RESET        : in    std_logic
); 
end component;

component FRAME_CHECK 
generic
(
    RX_DATA_WIDTH            : integer := 16;
    USE_COMMA                : integer := 1;
    NONE_MSB_FIRST_DEC       : integer := 0;
    CHANBOND_SEQ_LEN         : integer := 1;
    WORDS_IN_BRAM            : integer := 256;
    CONFIG_INDEPENDENT_LANES : integer := 0;
    START_OF_PACKET_CHAR     : std_logic_vector := x"55fb";
    MEM_00       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_01       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_02       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_03       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_04       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_05       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_06       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_07       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_08       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_09       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_0A       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_0B       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_0C       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_0D       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_0E       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_0F       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_10       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_11       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_12       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_13       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_14       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_15       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_16       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_17       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_18       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_19       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_1A       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_1B       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_1C       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_1D       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_1E       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_1F       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_20       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_21       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_22       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_23       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_24       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_25       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_26       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_27       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_28       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_29       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_2A       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_2B       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_2C       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_2D       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_2E       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_2F       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_30       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_31       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_32       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_33       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_34       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_35       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_36       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_37       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_38       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_39       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_3A       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_3B       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_3C       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_3D       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_3E       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_3F       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEMP_00      : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEMP_01      : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEMP_02      : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEMP_03      : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEMP_04      : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEMP_05      : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEMP_06      : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEMP_07      : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000"
);
port
(
    -- User Interface
    RX_DATA                  : in  std_logic_vector((RX_DATA_WIDTH-1) downto 0); 
    RX_ENMCOMMA_ALIGN        : out std_logic;
    RX_ENPCOMMA_ALIGN        : out std_logic;
    RX_ENCHAN_SYNC           : out std_logic; 
    RX_CHANBOND_SEQ          : in  std_logic; 

    -- Control Interface
    INC_IN                   : in std_logic; 
    INC_OUT                  : out std_logic; 
    PATTERN_MATCH_N          : out std_logic;
    RESET_ON_ERROR           : in std_logic; 
    
    -- Error Monitoring
    ERROR_COUNT              : out std_logic_vector(7 downto 0);

    -- Track Data
    TRACK_DATA               : out std_logic;

    -- System Interface
    USER_CLK                 : in std_logic;
    SYSTEM_RESET             : in std_logic
  
);
end component;

component MGT_USRCLK_SOURCE_PLL 
generic
(
    MULT                 : integer          := 2;
    DIVIDE               : integer          := 2;
    FEEDBACK             : string           := "CLKFBOUT";    
    CLK_PERIOD           : real             := 8.0;
    OUT0_DIVIDE          : integer          := 2;
    OUT1_DIVIDE          : integer          := 2;
    OUT2_DIVIDE          : integer          := 2;
    OUT3_DIVIDE          : integer          := 2   
);
port
( 
    CLK0_OUT                : out std_logic;
    CLK1_OUT                : out std_logic;
    CLK2_OUT                : out std_logic;
    CLK3_OUT                : out std_logic;
    CLK_IN                  : in  std_logic;
    CLKFB_IN                : in  std_logic;    
    CLKFB_OUT               : out std_logic;      
    PLL_LOCKED_OUT          : out std_logic;
    PLL_RESET_IN            : in  std_logic
);
end component;





-- Chipscope modules
attribute syn_black_box                : boolean;
attribute syn_noprune                  : boolean;


component shared_vio
port
(
    control                 : inout  std_logic_vector(35 downto 0);
    async_in                : in  std_logic_vector(31 downto 0);
    async_out               : out std_logic_vector(31 downto 0)
);
end component;
attribute syn_black_box of shared_vio : component is TRUE;
attribute syn_noprune of shared_vio   : component is TRUE;


component data_vio
port
(
    control                 : inout  std_logic_vector(35 downto 0);
    async_in                : in  std_logic_vector(139 downto 0);
    async_out               : out std_logic_vector(139 downto 0)
);
end component;
attribute syn_black_box of data_vio : component is TRUE;
attribute syn_noprune of data_vio   : component is TRUE;


component icon
port
(
    control0                : inout std_logic_vector(35 downto 0);
    control1                : inout std_logic_vector(35 downto 0);
    control2                : inout std_logic_vector(35 downto 0);
    control3                : inout std_logic_vector(35 downto 0);
    control4                : inout std_logic_vector(35 downto 0);
    control5                : inout std_logic_vector(35 downto 0);
    control6                : inout std_logic_vector(35 downto 0);
    control7                : inout std_logic_vector(35 downto 0);
    control8                : inout std_logic_vector(35 downto 0);
    control9                : inout std_logic_vector(35 downto 0);
    control10               : inout std_logic_vector(35 downto 0);
    control11               : inout std_logic_vector(35 downto 0);
    control12               : inout std_logic_vector(35 downto 0)
);
end component;
attribute syn_black_box of icon : component is TRUE;
attribute syn_noprune of icon   : component is TRUE;


component ila
port
(
    control                 : inout  std_logic_vector(35 downto 0);
    clk                     : in  std_logic;
    trig0                   : in  std_logic_vector(84 downto 0)
);
end component;
attribute syn_black_box of ila : component is TRUE;
attribute syn_noprune of ila   : component is TRUE;


component null_vio
port
(
    control                 : inout  std_logic_vector(35 downto 0)
);
end component;
attribute syn_black_box of null_vio : component is TRUE;
attribute syn_noprune of null_vio   : component is TRUE;


--***********************************Parameter Declarations********************

    constant DLY : time := 1 ns;
    
--************************** Register Declarations ****************************

    signal     tile0_tx_resetdone0_r           : std_logic;
    signal     tile0_tx_resetdone0_r2          : std_logic;
    signal     tile0_rx_resetdone0_r           : std_logic;
    signal     tile0_rx_resetdone0_r2          : std_logic;
    signal     tile0_tx_resetdone1_r           : std_logic;
    signal     tile0_tx_resetdone1_r2          : std_logic;
    signal     tile0_rx_resetdone1_r           : std_logic;
    signal     tile0_rx_resetdone1_r2          : std_logic;

--**************************** Wire Declarations ******************************

    -------------------------- MGT Wrapper Wires ------------------------------

    --________________________________________________________________________
    --________________________________________________________________________
    --TILE0   (X0_Y0)

    ------------------------ Loopback and Powerdown Ports ----------------------
    signal  tile0_loopback0_i               : std_logic_vector(2 downto 0);
    signal  tile0_loopback1_i               : std_logic_vector(2 downto 0);
    signal  tile0_rxpowerdown0_i            : std_logic_vector(1 downto 0);
    signal  tile0_rxpowerdown1_i            : std_logic_vector(1 downto 0);
    signal  tile0_txpowerdown0_i            : std_logic_vector(1 downto 0);
    signal  tile0_txpowerdown1_i            : std_logic_vector(1 downto 0);
    --------------------------------- PLL Ports --------------------------------
    signal  tile0_gtpreset0_i               : std_logic;
    signal  tile0_gtpreset1_i               : std_logic;
    signal  tile0_plllkdet0_i               : std_logic;
    signal  tile0_plllkdet1_i               : std_logic;
    signal  tile0_resetdone0_i              : std_logic;
    signal  tile0_resetdone1_i              : std_logic;
    ----------------------- Receive Ports - 8b10b Decoder ----------------------
    signal  tile0_rxchariscomma0_i          : std_logic;
    signal  tile0_rxchariscomma1_i          : std_logic;
    signal  tile0_rxcharisk0_i              : std_logic;
    signal  tile0_rxcharisk1_i              : std_logic;
    signal  tile0_rxdisperr0_i              : std_logic;
    signal  tile0_rxdisperr1_i              : std_logic;
    signal  tile0_rxnotintable0_i           : std_logic;
    signal  tile0_rxnotintable1_i           : std_logic;
    signal  tile0_rxrundisp0_i              : std_logic;
    signal  tile0_rxrundisp1_i              : std_logic;
    ---------------------- Receive Ports - Clock Correction --------------------
    signal  tile0_rxclkcorcnt0_i            : std_logic_vector(2 downto 0);
    signal  tile0_rxclkcorcnt1_i            : std_logic_vector(2 downto 0);
    --------------- Receive Ports - Comma Detection and Alignment --------------
    signal  tile0_rxenmcommaalign0_i        : std_logic;
    signal  tile0_rxenmcommaalign1_i        : std_logic;
    signal  tile0_rxenpcommaalign0_i        : std_logic;
    signal  tile0_rxenpcommaalign1_i        : std_logic;
    ------------------- Receive Ports - RX Data Path interface -----------------
    signal  tile0_rxdata0_i                 : std_logic_vector(7 downto 0);
    signal  tile0_rxdata1_i                 : std_logic_vector(7 downto 0);
    signal  tile0_rxrecclk0_i               : std_logic;
    signal  tile0_rxrecclk1_i               : std_logic;
    signal  tile0_rxreset0_i                : std_logic;
    signal  tile0_rxreset1_i                : std_logic;
    ----------- Receive Ports - RX Elastic Buffer and Phase Alignment ----------
    signal  tile0_rxbufreset0_i             : std_logic;
    signal  tile0_rxbufreset1_i             : std_logic;
    signal  tile0_rxbufstatus0_i            : std_logic_vector(2 downto 0);
    signal  tile0_rxbufstatus1_i            : std_logic_vector(2 downto 0);
    ---------------------------- TX/RX Datapath Ports --------------------------
    signal  tile0_gtpclkout0_i              : std_logic_vector(1 downto 0);
    signal  tile0_gtpclkout1_i              : std_logic_vector(1 downto 0);
    ------------------- Transmit Ports - 8b10b Encoder Control -----------------
    signal  tile0_txchardispmode0_i         : std_logic;
    signal  tile0_txchardispmode1_i         : std_logic;
    signal  tile0_txchardispval0_i          : std_logic;
    signal  tile0_txchardispval1_i          : std_logic;
    signal  tile0_txcharisk0_i              : std_logic;
    signal  tile0_txcharisk1_i              : std_logic;
    --------------- Transmit Ports - TX Buffer and Phase Alignment -------------
    signal  tile0_txbufstatus0_i            : std_logic_vector(1 downto 0);
    signal  tile0_txbufstatus1_i            : std_logic_vector(1 downto 0);
    ------------------ Transmit Ports - TX Data Path interface -----------------
    signal  tile0_txdata0_i                 : std_logic_vector(7 downto 0);
    signal  tile0_txdata1_i                 : std_logic_vector(7 downto 0);
    signal  tile0_txoutclk0_i               : std_logic;
    signal  tile0_txoutclk1_i               : std_logic;
    signal  tile0_txreset0_i                : std_logic;
    signal  tile0_txreset1_i                : std_logic;


    ------------------------------- Global Signals -----------------------------
    signal  tile0_tx_system_reset0_c        : std_logic;
    signal  tile0_rx_system_reset0_c        : std_logic;
    signal  tile0_tx_system_reset1_c        : std_logic;
    signal  tile0_rx_system_reset1_c        : std_logic;
    signal  tied_to_ground_i                : std_logic;
    signal  tied_to_ground_vec_i            : std_logic_vector(191 downto 0);
    signal  tied_to_vcc_i                   : std_logic;
    signal  tied_to_vcc_vec_i               : std_logic_vector(7 downto 0);
    signal  drp_clk_in_i                    : std_logic;
    signal  tile0_refclkout_bufg_i          : std_logic;
    
    
    ----------------------------- User Clocks ---------------------------------
    signal  tile0_txusrclk0_i               : std_logic;
    signal  tile0_gtpclkout0_0_to_bufg_i    : std_logic;


    ----------------------- Frame check/gen Module Signals --------------------
    signal  tile0_gtp0_refclk_i             : std_logic;
    signal  tile0_matchn0_i                 : std_logic;
    
    signal  tile0_txcharisk0_float_i        : std_logic_vector(2 downto 0);
    signal  tile0_txdata0_float_i           : std_logic_vector(31 downto 0);
    signal  tile0_track_data0_i             : std_logic;
    signal  tile0_error_count0_i            : std_logic_vector(7 downto 0);
    signal  tile0_frame_check0_reset_i      : std_logic;
    signal  tile0_inc_in0_i                 : std_logic;
    signal  tile0_inc_out0_i                : std_logic;
    signal  tile0_matchn1_i                 : std_logic;
    
    signal  tile0_txcharisk1_float_i        : std_logic_vector(2 downto 0);
    signal  tile0_txdata1_float_i           : std_logic_vector(31 downto 0);
    signal  tile0_track_data1_i             : std_logic;
    signal  tile0_error_count1_i            : std_logic_vector(7 downto 0);
    signal  tile0_frame_check1_reset_i      : std_logic;
    signal  tile0_inc_in1_i                 : std_logic;
    signal  tile0_inc_out1_i                : std_logic;

    signal  reset_on_data_error_i           : std_logic;
    signal  track_data_out_i                : std_logic;
    
    ------------------------- Sync Module Signals -----------------------------

    ----------------------- Chipscope Signals ---------------------------------

    signal  shared_vio_control_i            : std_logic_vector(35 downto 0);
    signal  tile0_data_vio_control_i        : std_logic_vector(35 downto 0);
    signal  tile0_gtp0_ila_control_i        : std_logic_vector(35 downto 0);
    signal  tile0_gtp1_ila_control_i        : std_logic_vector(35 downto 0);
    signal  null_vio_4_i                    : std_logic_vector(35 downto 0);
    signal  null_vio_5_i                    : std_logic_vector(35 downto 0);
    signal  null_vio_6_i                    : std_logic_vector(35 downto 0);
    signal  null_vio_7_i                    : std_logic_vector(35 downto 0);
    signal  null_vio_8_i                    : std_logic_vector(35 downto 0);
    signal  null_vio_9_i                    : std_logic_vector(35 downto 0);
    signal  null_vio_10_i                   : std_logic_vector(35 downto 0);
    signal  null_vio_11_i                   : std_logic_vector(35 downto 0);
    signal  null_vio_12_i                   : std_logic_vector(35 downto 0);
    signal  shared_vio_in_i                 : std_logic_vector(31 downto 0);
    signal  shared_vio_out_i                : std_logic_vector(31 downto 0);

    signal  tile0_data_vio_in_i             : std_logic_vector(139 downto 0);
    signal  tile0_data_vio_out_i            : std_logic_vector(139 downto 0);
    signal  tile0_ila_in0_i                 : std_logic_vector(84 downto 0);
    signal  tile0_ila_in1_i                 : std_logic_vector(84 downto 0);


    signal  gtpreset0_i                     : std_logic;
    signal  gtpreset1_i                     : std_logic;
    signal  user_tx_reset_i                 : std_logic;
    signal  user_rx_reset_i                 : std_logic;

--**************************** Main Body of Code *******************************
begin

    --  Static signal Assigments
    tied_to_ground_i                        <= '0';
    tied_to_ground_vec_i                    <= x"000000000000000000000000000000000000000000000000";
    tied_to_vcc_i                           <= '1';
    tied_to_vcc_vec_i                       <= x"ff";


    


    -----------------------Dedicated GTP Reference Clock Inputs ---------------
    -- The dedicated reference clock inputs you selected in the GUI are implemented using
    -- IBUFDS instances.
    --
    -- In the UCF file for this example design, you will see that each of
    -- these IBUFDS instances has been LOCed to a particular set of pins. By LOCing to these
    -- locations, we tell the tools to use the dedicated input buffers to the GTP reference
    -- clock network, rather than general purpose IOs. To select other pins, consult the 
    -- Implementation chapter of UG___, or rerun the wizard.
    --
    -- This network is the highest performace (lowest jitter) option for providing clocks
    -- to the GTP transceivers.
    
    tile0_gtp0_refclk_ibufds_i : IBUFDS
    port map
    (
        O                               =>      tile0_gtp0_refclk_i,
        I                               =>      tile0_gtp0_REFCLK_PAD_P_IN,
        IB                              =>      tile0_gtp0_REFCLK_PAD_N_IN
    );

    ----------------------------------- User Clocks ---------------------------
    
    -- The clock resources in this section were added based on userclk source selections on
    -- the Latency, Buffering, and Clocking page of the GUI. A few notes about user clocks:
    -- * The userclk and userclk2 for each GTP datapath (TX and RX) must be phase aligned to 
    --   avoid data errors in the fabric interface whenever the datapath is wider than 10 bits
    -- * To minimize clock resources, you can share clocks between GTPs. GTPs using the same frequency
    --   or multiples of the same frequency can be accomadated using DCMs and PLLs. Use caution when
    --   using RXRECCLK as a clock source, however - these clocks can typically only be shared if all
    --   the channels using the clock are receiving data from TX channels that share a reference clock 
    --   source with each other.

    gtpclkout0_0_bufg0_bufio2_i : BUFIO2
    generic map
    (
        DIVIDE                          =>      1,
        DIVIDE_BYPASS                   =>      TRUE
    )
    port map
    (
        I                               =>      tile0_gtpclkout0_i(0),
        DIVCLK                          =>      tile0_gtpclkout0_0_to_bufg_i,
        IOCLK                           =>      open,
        SERDESSTROBE                    =>      open
    );

    gtpclkout0_0_bufg0_i : BUFG
    port map
    (
        I                               =>      tile0_gtpclkout0_0_to_bufg_i,
        O                               =>      tile0_txusrclk0_i
    );






    ----------------------------- The GTP Wrapper -----------------------------
    
    -- Use the instantiation template in the top directory to add the GTP wrapper to your design.
    -- In this example, the wrapper is wired up for basic operation with a frame generator and frame 
    -- checker. The GTPs will reset, then attempt to align and transmit data. If channel bonding is 
    -- enabled, bonding should occur after alignment.
    

    -- Wire all PLLLKDET signals to the top level as output ports
    TILE0_GTP0_PLLLKDET_OUT                 <= tile0_plllkdet0_i;

    -- Hold the TX in reset till the TX user clocks are stable
    tile0_txreset0_i                    <= not tile0_plllkdet0_i;
    tile0_txreset1_i                    <= not tile0_plllkdet0_i;

    -- Hold the RX in reset till the RX user clocks are stable
    tile0_rxreset0_i                    <= not tile0_plllkdet0_i;
    tile0_rxreset1_i                    <= not tile0_plllkdet0_i;

    pcs_pma_s6_gtpwizard_i : pcs_pma_s6_gtpwizard
    generic map
    (
        WRAPPER_SIM_GTPRESET_SPEEDUP    =>      EXAMPLE_SIM_GTPRESET_SPEEDUP,
        WRAPPER_CLK25_DIVIDER_0         =>      5,
        WRAPPER_CLK25_DIVIDER_1         =>      5,
        WRAPPER_PLL_DIVSEL_FB_0         =>      2,
        WRAPPER_PLL_DIVSEL_FB_1         =>      2,
        WRAPPER_PLL_DIVSEL_REF_0        =>      1,
        WRAPPER_PLL_DIVSEL_REF_1        =>      1,
        WRAPPER_SIMULATION              =>      EXAMPLE_SIMULATION
    )
    port map
    (
 
 
 
 
 
        --_____________________________________________________________________
        --_____________________________________________________________________
        --TILE0  (X0_Y0)

        ------------------------ Loopback and Powerdown Ports ----------------------
        TILE0_LOOPBACK0_IN              =>      tile0_loopback0_i,
        TILE0_LOOPBACK1_IN              =>      tile0_loopback1_i,
        TILE0_RXPOWERDOWN0_IN           =>      tile0_rxpowerdown0_i,
        TILE0_RXPOWERDOWN1_IN           =>      tile0_rxpowerdown1_i,
        TILE0_TXPOWERDOWN0_IN           =>      tile0_txpowerdown0_i,
        TILE0_TXPOWERDOWN1_IN           =>      tile0_txpowerdown1_i,
        --------------------------------- PLL Ports --------------------------------
        TILE0_CLK00_IN                  =>      tile0_gtp0_refclk_i,
        TILE0_CLK01_IN                  =>      tied_to_ground_i,
        TILE0_GTPRESET0_IN              =>      tile0_gtpreset0_i,
        TILE0_GTPRESET1_IN              =>      tile0_gtpreset0_i,
        TILE0_PLLLKDET0_OUT             =>      tile0_plllkdet0_i,
        TILE0_RESETDONE0_OUT            =>      tile0_resetdone0_i,
        TILE0_RESETDONE1_OUT            =>      tile0_resetdone1_i,
        ----------------------- Receive Ports - 8b10b Decoder ----------------------
        TILE0_RXCHARISCOMMA0_OUT        =>      tile0_rxchariscomma0_i,
        TILE0_RXCHARISCOMMA1_OUT        =>      tile0_rxchariscomma1_i,
        TILE0_RXCHARISK0_OUT            =>      tile0_rxcharisk0_i,
        TILE0_RXCHARISK1_OUT            =>      tile0_rxcharisk1_i,
        TILE0_RXDISPERR0_OUT            =>      tile0_rxdisperr0_i,
        TILE0_RXDISPERR1_OUT            =>      tile0_rxdisperr1_i,
        TILE0_RXNOTINTABLE0_OUT         =>      tile0_rxnotintable0_i,
        TILE0_RXNOTINTABLE1_OUT         =>      tile0_rxnotintable1_i,
        TILE0_RXRUNDISP0_OUT            =>      tile0_rxrundisp0_i,
        TILE0_RXRUNDISP1_OUT            =>      tile0_rxrundisp1_i,
        ---------------------- Receive Ports - Clock Correction --------------------
        TILE0_RXCLKCORCNT0_OUT          =>      tile0_rxclkcorcnt0_i,
        TILE0_RXCLKCORCNT1_OUT          =>      tile0_rxclkcorcnt1_i,
        --------------- Receive Ports - Comma Detection and Alignment --------------
        TILE0_RXENMCOMMAALIGN0_IN       =>      tile0_rxenmcommaalign0_i,
        TILE0_RXENMCOMMAALIGN1_IN       =>      tile0_rxenmcommaalign1_i,
        TILE0_RXENPCOMMAALIGN0_IN       =>      tile0_rxenpcommaalign0_i,
        TILE0_RXENPCOMMAALIGN1_IN       =>      tile0_rxenpcommaalign1_i,
        ------------------- Receive Ports - RX Data Path interface -----------------
        TILE0_RXDATA0_OUT               =>      tile0_rxdata0_i,
        TILE0_RXDATA1_OUT               =>      tile0_rxdata1_i,
        TILE0_RXRECCLK0_OUT             =>      tile0_rxrecclk0_i,
        TILE0_RXRECCLK1_OUT             =>      tile0_rxrecclk1_i,
        TILE0_RXRESET0_IN               =>      tile0_rxreset0_i,
        TILE0_RXRESET1_IN               =>      tile0_rxreset1_i,
        TILE0_RXUSRCLK0_IN              =>      tile0_txusrclk0_i,
        TILE0_RXUSRCLK1_IN              =>      tile0_txusrclk0_i,
        TILE0_RXUSRCLK20_IN             =>      tile0_txusrclk0_i,
        TILE0_RXUSRCLK21_IN             =>      tile0_txusrclk0_i,
        ------- Receive Ports - RX Driver,OOB signalling,Coupling and Eq.,CDR ------
        TILE0_RXN0_IN                   =>      RXN_IN(0),
        TILE0_RXN1_IN                   =>      RXN_IN(1),
        TILE0_RXP0_IN                   =>      RXP_IN(0),
        TILE0_RXP1_IN                   =>      RXP_IN(1),
        ----------- Receive Ports - RX Elastic Buffer and Phase Alignment ----------
        TILE0_RXBUFRESET0_IN            =>      tile0_rxbufreset0_i,
        TILE0_RXBUFRESET1_IN            =>      tile0_rxbufreset1_i,
        TILE0_RXBUFSTATUS0_OUT          =>      tile0_rxbufstatus0_i,
        TILE0_RXBUFSTATUS1_OUT          =>      tile0_rxbufstatus1_i,
        ---------------------------- TX/RX Datapath Ports --------------------------
        TILE0_GTPCLKOUT0_OUT            =>      tile0_gtpclkout0_i,
        TILE0_GTPCLKOUT1_OUT            =>      tile0_gtpclkout1_i,
        ------------------- Transmit Ports - 8b10b Encoder Control -----------------
        TILE0_TXCHARDISPMODE0_IN        =>      tile0_txchardispmode0_i,
        TILE0_TXCHARDISPMODE1_IN        =>      tile0_txchardispmode1_i,
        TILE0_TXCHARDISPVAL0_IN         =>      tile0_txchardispval0_i,
        TILE0_TXCHARDISPVAL1_IN         =>      tile0_txchardispval1_i,
        TILE0_TXCHARISK0_IN             =>      tile0_txcharisk0_i,
        TILE0_TXCHARISK1_IN             =>      tile0_txcharisk1_i,
        --------------- Transmit Ports - TX Buffer and Phase Alignment -------------
        TILE0_TXBUFSTATUS0_OUT          =>      tile0_txbufstatus0_i,
        TILE0_TXBUFSTATUS1_OUT          =>      tile0_txbufstatus1_i,
        ------------------ Transmit Ports - TX Data Path interface -----------------
        TILE0_TXDATA0_IN                =>      tile0_txdata0_i,
        TILE0_TXDATA1_IN                =>      tile0_txdata1_i,
        TILE0_TXOUTCLK0_OUT             =>      tile0_txoutclk0_i,
        TILE0_TXOUTCLK1_OUT             =>      tile0_txoutclk1_i,
        TILE0_TXRESET0_IN               =>      tile0_txreset0_i,
        TILE0_TXRESET1_IN               =>      tile0_txreset1_i,
        TILE0_TXUSRCLK0_IN              =>      tile0_txusrclk0_i,
        TILE0_TXUSRCLK1_IN              =>      tile0_txusrclk0_i,
        TILE0_TXUSRCLK20_IN             =>      tile0_txusrclk0_i,
        TILE0_TXUSRCLK21_IN             =>      tile0_txusrclk0_i,
        --------------- Transmit Ports - TX Driver and OOB signalling --------------
        TILE0_TXN0_OUT                  =>      TXN_OUT(0),
        TILE0_TXN1_OUT                  =>      TXN_OUT(1),
        TILE0_TXP0_OUT                  =>      TXP_OUT(0),
        TILE0_TXP1_OUT                  =>      TXP_OUT(1)


    );







    -------------------------- User Module Resets -----------------------------
    -- All the User Modules i.e. FRAME_GEN, FRAME_CHECK and the sync modules
    -- are held in reset till the RESETDONE goes high. 
    -- The RESETDONE is registered a couple of times on USRCLK2 and connected 
    -- to the reset of the modules
    
    process( tile0_txusrclk0_i,tile0_resetdone0_i)
    begin
        if(tile0_resetdone0_i = '0') then
            tile0_rx_resetdone0_r  <= '0'   ;
            tile0_rx_resetdone0_r2 <= '0'   ;
        elsif(tile0_txusrclk0_i'event and tile0_txusrclk0_i = '1') then
            tile0_rx_resetdone0_r  <= tile0_resetdone0_i   ;
            tile0_rx_resetdone0_r2 <= tile0_rx_resetdone0_r   ;
        end if;
    end process;
    
    process( tile0_txusrclk0_i,tile0_resetdone1_i)
    begin
        if(tile0_resetdone1_i = '0') then
            tile0_rx_resetdone1_r  <= '0'   ;
            tile0_rx_resetdone1_r2 <= '0'   ;
        elsif(tile0_txusrclk0_i'event and tile0_txusrclk0_i = '1') then
            tile0_rx_resetdone1_r  <= tile0_resetdone1_i   ;
            tile0_rx_resetdone1_r2 <= tile0_rx_resetdone1_r   ;
        end if;
    end process;
    
    process( tile0_txusrclk0_i,tile0_resetdone0_i)
    begin
        if (tile0_resetdone0_i = '0') then 
            tile0_tx_resetdone0_r    <=   '0'   ;
            tile0_tx_resetdone0_r2   <=   '0'   ;
        elsif(tile0_txusrclk0_i'event and tile0_txusrclk0_i = '1') then
            tile0_tx_resetdone0_r    <=   tile0_resetdone0_i  ;
            tile0_tx_resetdone0_r2   <=   tile0_tx_resetdone0_r   ;
        end if;
    end process; 
    process( tile0_txusrclk0_i,tile0_resetdone1_i)
    begin
        if (tile0_resetdone1_i = '0') then 
            tile0_tx_resetdone1_r    <=   '0'   ;
            tile0_tx_resetdone1_r2   <=   '0'   ;
        elsif(tile0_txusrclk0_i'event and tile0_txusrclk0_i = '1') then
            tile0_tx_resetdone1_r    <=   tile0_resetdone1_i  ;
            tile0_tx_resetdone1_r2   <=   tile0_tx_resetdone1_r   ;
        end if;
    end process; 

    ------------------------------ Frame Generators ---------------------------
    -- The example design uses Block RAM based frame generators to provide test
    -- data to the GTPs for transmission. By default the frame generators are 
    -- loaded with an incrementing data sequence that includes commas/alignment
    -- characters for alignment. If your protocol uses channel bonding, the 
    -- frame generator will also be preloaded with a channel bonding sequence.
    
    -- You can modify the data transmitted by changing the INIT values of the frame
    -- generator in this file. Pay careful attention to bit order and the spacing
    -- of your control and alignment characters.

    tile0_frame_gen0 : FRAME_GEN
    generic map
    (
        WORDS_IN_BRAM                   =>      EXAMPLE_WORDS_IN_BRAM,
        MEM_00                  =>  x"0000000600000005000000040000000300000002000000bc0000000100000000",
        MEM_01                  =>  x"0000000e0000000d0000000c0000000b0000000a000000090000000800000007",
        MEM_02                  =>  x"000000160000001500000014000000130000001200000011000000100000000f",
        MEM_03                  =>  x"0000001e0000001d0000001c0000001b0000001a000000190000001800000017",
        MEM_04                  =>  x"000000260000002500000024000000230000002200000021000000200000001f",
        MEM_05                  =>  x"0000002e0000002d0000002c0000002b0000002a000000290000002800000027",
        MEM_06                  =>  x"000000360000003500000034000000330000003200000031000000300000002f",
        MEM_07                  =>  x"0000003e0000003d0000003c0000003b0000003a000000390000003800000037",
        MEM_08                  =>  x"000000460000004500000044000000430000004200000041000000400000003f",
        MEM_09                  =>  x"0000004e0000004d0000004c0000004b0000004a000000490000004800000047",
        MEM_0A                  =>  x"000000560000005500000054000000530000005200000051000000500000004f",
        MEM_0B                  =>  x"0000005e0000005d0000005c0000005b0000005a000000590000005800000057",
        MEM_0C                  =>  x"000000660000006500000064000000630000006200000061000000600000005f",
        MEM_0D                  =>  x"0000006e0000006d0000006c0000006b0000006a000000690000006800000067",
        MEM_0E                  =>  x"000000760000007500000074000000730000007200000071000000700000006f",
        MEM_0F                  =>  x"0000007e0000007d0000007c0000007b0000007a000000790000007800000077",
        MEM_10                  =>  x"0000000600000005000000040000000300000002000000bc0000000100000000",
        MEM_11                  =>  x"0000000e0000000d0000000c0000000b0000000a000000090000000800000007",
        MEM_12                  =>  x"000000160000001500000014000000130000001200000011000000100000000f",
        MEM_13                  =>  x"0000001e0000001d0000001c0000001b0000001a000000190000001800000017",
        MEM_14                  =>  x"000000260000002500000024000000230000002200000021000000200000001f",
        MEM_15                  =>  x"0000002e0000002d0000002c0000002b0000002a000000290000002800000027",
        MEM_16                  =>  x"000000360000003500000034000000330000003200000031000000300000002f",
        MEM_17                  =>  x"0000003e0000003d0000003c0000003b0000003a000000390000003800000037",
        MEM_18                  =>  x"000000460000004500000044000000430000004200000041000000400000003f",
        MEM_19                  =>  x"0000004e0000004d0000004c0000004b0000004a000000490000004800000047",
        MEM_1A                  =>  x"000000560000005500000054000000530000005200000051000000500000004f",
        MEM_1B                  =>  x"0000005e0000005d0000005c0000005b0000005a000000590000005800000057",
        MEM_1C                  =>  x"000000660000006500000064000000630000006200000061000000600000005f",
        MEM_1D                  =>  x"0000006e0000006d0000006c0000006b0000006a000000690000006800000067",
        MEM_1E                  =>  x"000000760000007500000074000000730000007200000071000000700000006f",
        MEM_1F                  =>  x"0000007e0000007d0000007c0000007b0000007a000000790000007800000077",
        MEM_20                  =>  x"0000000600000005000000040000000300000002000000bc0000000100000000",
        MEM_21                  =>  x"0000000e0000000d0000000c0000000b0000000a000000090000000800000007",
        MEM_22                  =>  x"000000160000001500000014000000130000001200000011000000100000000f",
        MEM_23                  =>  x"0000001e0000001d0000001c0000001b0000001a000000190000001800000017",
        MEM_24                  =>  x"000000260000002500000024000000230000002200000021000000200000001f",
        MEM_25                  =>  x"0000002e0000002d0000002c0000002b0000002a000000290000002800000027",
        MEM_26                  =>  x"000000360000003500000034000000330000003200000031000000300000002f",
        MEM_27                  =>  x"0000003e0000003d0000003c0000003b0000003a000000390000003800000037",
        MEM_28                  =>  x"000000460000004500000044000000430000004200000041000000400000003f",
        MEM_29                  =>  x"0000004e0000004d0000004c0000004b0000004a000000490000004800000047",
        MEM_2A                  =>  x"000000560000005500000054000000530000005200000051000000500000004f",
        MEM_2B                  =>  x"0000005e0000005d0000005c0000005b0000005a000000590000005800000057",
        MEM_2C                  =>  x"000000660000006500000064000000630000006200000061000000600000005f",
        MEM_2D                  =>  x"0000006e0000006d0000006c0000006b0000006a000000690000006800000067",
        MEM_2E                  =>  x"000000760000007500000074000000730000007200000071000000700000006f",
        MEM_2F                  =>  x"0000007e0000007d0000007c0000007b0000007a000000790000007800000077",
        MEM_30                  =>  x"0000000600000005000000040000000300000002000000bc0000000100000000",
        MEM_31                  =>  x"0000000e0000000d0000000c0000000b0000000a000000090000000800000007",
        MEM_32                  =>  x"000000160000001500000014000000130000001200000011000000100000000f",
        MEM_33                  =>  x"0000001e0000001d0000001c0000001b0000001a000000190000001800000017",
        MEM_34                  =>  x"000000260000002500000024000000230000002200000021000000200000001f",
        MEM_35                  =>  x"0000002e0000002d0000002c0000002b0000002a000000290000002800000027",
        MEM_36                  =>  x"000000360000003500000034000000330000003200000031000000300000002f",
        MEM_37                  =>  x"0000003e0000003d0000003c0000003b0000003a000000390000003800000037",
        MEM_38                  =>  x"000000460000004500000044000000430000004200000041000000400000003f",
        MEM_39                  =>  x"0000004e0000004d0000004c0000004b0000004a000000490000004800000047",
        MEM_3A                  =>  x"000000560000005500000054000000530000005200000051000000500000004f",
        MEM_3B                  =>  x"0000005e0000005d0000005c0000005b0000005a000000590000005800000057",
        MEM_3C                  =>  x"000000660000006500000064000000630000006200000061000000600000005f",
        MEM_3D                  =>  x"0000006e0000006d0000006c0000006b0000006a000000690000006800000067",
        MEM_3E                  =>  x"000000760000007500000074000000730000007200000071000000700000006f",
        MEM_3F                  =>  x"0000007e0000007d0000007c0000007b0000007a000000790000007800000077",
        MEMP_00                  =>  x"0000000000000000000000000000000000000000000000000000000000000100",
        MEMP_01                  =>  x"0000000000000000000000000000000000000000000000000000000000000000",
        MEMP_02                  =>  x"0000000000000000000000000000000000000000000000000000000000000100",
        MEMP_03                  =>  x"0000000000000000000000000000000000000000000000000000000000000000",
        MEMP_04                  =>  x"0000000000000000000000000000000000000000000000000000000000000100",
        MEMP_05                  =>  x"0000000000000000000000000000000000000000000000000000000000000000",
        MEMP_06                  =>  x"0000000000000000000000000000000000000000000000000000000000000100",
        MEMP_07                  =>  x"0000000000000000000000000000000000000000000000000000000000000000"
    )
    port map
    (
        -- User Interface
        TX_DATA(39 downto 8)            =>      tile0_txdata0_float_i,
        TX_DATA(7 downto 0)             =>      tile0_txdata0_i,
 
        TX_CHARISK(3 downto 1)          =>      tile0_txcharisk0_float_i,
        TX_CHARISK(0)                   =>      tile0_txcharisk0_i,
        -- System Interface
        USER_CLK                        =>      tile0_txusrclk0_i,
        SYSTEM_RESET                    =>      tile0_tx_system_reset0_c
    );
    
    tile0_frame_gen1 : FRAME_GEN
    generic map
    (
        WORDS_IN_BRAM                   =>      EXAMPLE_WORDS_IN_BRAM,
        MEM_00                  =>  x"0000000600000005000000040000000300000002000000bc0000000100000000",
        MEM_01                  =>  x"0000000e0000000d0000000c0000000b0000000a000000090000000800000007",
        MEM_02                  =>  x"000000160000001500000014000000130000001200000011000000100000000f",
        MEM_03                  =>  x"0000001e0000001d0000001c0000001b0000001a000000190000001800000017",
        MEM_04                  =>  x"000000260000002500000024000000230000002200000021000000200000001f",
        MEM_05                  =>  x"0000002e0000002d0000002c0000002b0000002a000000290000002800000027",
        MEM_06                  =>  x"000000360000003500000034000000330000003200000031000000300000002f",
        MEM_07                  =>  x"0000003e0000003d0000003c0000003b0000003a000000390000003800000037",
        MEM_08                  =>  x"000000460000004500000044000000430000004200000041000000400000003f",
        MEM_09                  =>  x"0000004e0000004d0000004c0000004b0000004a000000490000004800000047",
        MEM_0A                  =>  x"000000560000005500000054000000530000005200000051000000500000004f",
        MEM_0B                  =>  x"0000005e0000005d0000005c0000005b0000005a000000590000005800000057",
        MEM_0C                  =>  x"000000660000006500000064000000630000006200000061000000600000005f",
        MEM_0D                  =>  x"0000006e0000006d0000006c0000006b0000006a000000690000006800000067",
        MEM_0E                  =>  x"000000760000007500000074000000730000007200000071000000700000006f",
        MEM_0F                  =>  x"0000007e0000007d0000007c0000007b0000007a000000790000007800000077",
        MEM_10                  =>  x"0000000600000005000000040000000300000002000000bc0000000100000000",
        MEM_11                  =>  x"0000000e0000000d0000000c0000000b0000000a000000090000000800000007",
        MEM_12                  =>  x"000000160000001500000014000000130000001200000011000000100000000f",
        MEM_13                  =>  x"0000001e0000001d0000001c0000001b0000001a000000190000001800000017",
        MEM_14                  =>  x"000000260000002500000024000000230000002200000021000000200000001f",
        MEM_15                  =>  x"0000002e0000002d0000002c0000002b0000002a000000290000002800000027",
        MEM_16                  =>  x"000000360000003500000034000000330000003200000031000000300000002f",
        MEM_17                  =>  x"0000003e0000003d0000003c0000003b0000003a000000390000003800000037",
        MEM_18                  =>  x"000000460000004500000044000000430000004200000041000000400000003f",
        MEM_19                  =>  x"0000004e0000004d0000004c0000004b0000004a000000490000004800000047",
        MEM_1A                  =>  x"000000560000005500000054000000530000005200000051000000500000004f",
        MEM_1B                  =>  x"0000005e0000005d0000005c0000005b0000005a000000590000005800000057",
        MEM_1C                  =>  x"000000660000006500000064000000630000006200000061000000600000005f",
        MEM_1D                  =>  x"0000006e0000006d0000006c0000006b0000006a000000690000006800000067",
        MEM_1E                  =>  x"000000760000007500000074000000730000007200000071000000700000006f",
        MEM_1F                  =>  x"0000007e0000007d0000007c0000007b0000007a000000790000007800000077",
        MEM_20                  =>  x"0000000600000005000000040000000300000002000000bc0000000100000000",
        MEM_21                  =>  x"0000000e0000000d0000000c0000000b0000000a000000090000000800000007",
        MEM_22                  =>  x"000000160000001500000014000000130000001200000011000000100000000f",
        MEM_23                  =>  x"0000001e0000001d0000001c0000001b0000001a000000190000001800000017",
        MEM_24                  =>  x"000000260000002500000024000000230000002200000021000000200000001f",
        MEM_25                  =>  x"0000002e0000002d0000002c0000002b0000002a000000290000002800000027",
        MEM_26                  =>  x"000000360000003500000034000000330000003200000031000000300000002f",
        MEM_27                  =>  x"0000003e0000003d0000003c0000003b0000003a000000390000003800000037",
        MEM_28                  =>  x"000000460000004500000044000000430000004200000041000000400000003f",
        MEM_29                  =>  x"0000004e0000004d0000004c0000004b0000004a000000490000004800000047",
        MEM_2A                  =>  x"000000560000005500000054000000530000005200000051000000500000004f",
        MEM_2B                  =>  x"0000005e0000005d0000005c0000005b0000005a000000590000005800000057",
        MEM_2C                  =>  x"000000660000006500000064000000630000006200000061000000600000005f",
        MEM_2D                  =>  x"0000006e0000006d0000006c0000006b0000006a000000690000006800000067",
        MEM_2E                  =>  x"000000760000007500000074000000730000007200000071000000700000006f",
        MEM_2F                  =>  x"0000007e0000007d0000007c0000007b0000007a000000790000007800000077",
        MEM_30                  =>  x"0000000600000005000000040000000300000002000000bc0000000100000000",
        MEM_31                  =>  x"0000000e0000000d0000000c0000000b0000000a000000090000000800000007",
        MEM_32                  =>  x"000000160000001500000014000000130000001200000011000000100000000f",
        MEM_33                  =>  x"0000001e0000001d0000001c0000001b0000001a000000190000001800000017",
        MEM_34                  =>  x"000000260000002500000024000000230000002200000021000000200000001f",
        MEM_35                  =>  x"0000002e0000002d0000002c0000002b0000002a000000290000002800000027",
        MEM_36                  =>  x"000000360000003500000034000000330000003200000031000000300000002f",
        MEM_37                  =>  x"0000003e0000003d0000003c0000003b0000003a000000390000003800000037",
        MEM_38                  =>  x"000000460000004500000044000000430000004200000041000000400000003f",
        MEM_39                  =>  x"0000004e0000004d0000004c0000004b0000004a000000490000004800000047",
        MEM_3A                  =>  x"000000560000005500000054000000530000005200000051000000500000004f",
        MEM_3B                  =>  x"0000005e0000005d0000005c0000005b0000005a000000590000005800000057",
        MEM_3C                  =>  x"000000660000006500000064000000630000006200000061000000600000005f",
        MEM_3D                  =>  x"0000006e0000006d0000006c0000006b0000006a000000690000006800000067",
        MEM_3E                  =>  x"000000760000007500000074000000730000007200000071000000700000006f",
        MEM_3F                  =>  x"0000007e0000007d0000007c0000007b0000007a000000790000007800000077",
        MEMP_00                  =>  x"0000000000000000000000000000000000000000000000000000000000000100",
        MEMP_01                  =>  x"0000000000000000000000000000000000000000000000000000000000000000",
        MEMP_02                  =>  x"0000000000000000000000000000000000000000000000000000000000000100",
        MEMP_03                  =>  x"0000000000000000000000000000000000000000000000000000000000000000",
        MEMP_04                  =>  x"0000000000000000000000000000000000000000000000000000000000000100",
        MEMP_05                  =>  x"0000000000000000000000000000000000000000000000000000000000000000",
        MEMP_06                  =>  x"0000000000000000000000000000000000000000000000000000000000000100",
        MEMP_07                  =>  x"0000000000000000000000000000000000000000000000000000000000000000"
    )
    port map
    (
        -- User Interface
        TX_DATA(39 downto 8)            =>      tile0_txdata1_float_i,
        TX_DATA(7 downto 0)             =>      tile0_txdata1_i,
 
        TX_CHARISK(3 downto 1)          =>      tile0_txcharisk1_float_i,
        TX_CHARISK(0)                   =>      tile0_txcharisk1_i,
        -- System Interface
        USER_CLK                        =>      tile0_txusrclk0_i,
        SYSTEM_RESET                    =>      tile0_tx_system_reset1_c
    );
    


    ---------------------------------- Frame Checkers -------------------------
    -- The example design uses Block RAM based frame checkers to verify incoming  
    -- data. By default the frame generators are loaded with a data sequence that 
    -- matches the outgoing sequence of the frame generators for the TX ports.
    
    -- You can modify the expected data sequence by changing the INIT values of the frame
    -- checkers in this file. Pay careful attention to bit order and the spacing
    -- of your control and alignment characters.
    
    -- When the frame checker receives data, it attempts to synchronise to the 
    -- incoming pattern by looking for the first sequence in the pattern. Once it 
    -- finds the first sequence, it increments through the sequence, and indicates an 
    -- error whenever the next value received does not match the expected value.

    tile0_frame_check0_reset_i              <= reset_on_data_error_i when (EXAMPLE_CONFIG_INDEPENDENT_LANES=0) else tile0_matchn0_i;

    -- tile0_frame_check0 is always connected to the lane with the start of char
    -- and this lane starts off the data checking on all the other lanes. The INC_IN port is tied off
    tile0_inc_in0_i                         <= '0';

    tile0_frame_check0 : FRAME_CHECK
    generic map
    (
        RX_DATA_WIDTH                   =>      8,
        USE_COMMA                       =>      1,
        WORDS_IN_BRAM                   =>      EXAMPLE_WORDS_IN_BRAM,
        CONFIG_INDEPENDENT_LANES        =>      1,
        START_OF_PACKET_CHAR            =>      x"bc",
        MEM_00                  =>  x"0000000600000005000000040000000300000002000000bc0000000100000000",
        MEM_01                  =>  x"0000000e0000000d0000000c0000000b0000000a000000090000000800000007",
        MEM_02                  =>  x"000000160000001500000014000000130000001200000011000000100000000f",
        MEM_03                  =>  x"0000001e0000001d0000001c0000001b0000001a000000190000001800000017",
        MEM_04                  =>  x"000000260000002500000024000000230000002200000021000000200000001f",
        MEM_05                  =>  x"0000002e0000002d0000002c0000002b0000002a000000290000002800000027",
        MEM_06                  =>  x"000000360000003500000034000000330000003200000031000000300000002f",
        MEM_07                  =>  x"0000003e0000003d0000003c0000003b0000003a000000390000003800000037",
        MEM_08                  =>  x"000000460000004500000044000000430000004200000041000000400000003f",
        MEM_09                  =>  x"0000004e0000004d0000004c0000004b0000004a000000490000004800000047",
        MEM_0A                  =>  x"000000560000005500000054000000530000005200000051000000500000004f",
        MEM_0B                  =>  x"0000005e0000005d0000005c0000005b0000005a000000590000005800000057",
        MEM_0C                  =>  x"000000660000006500000064000000630000006200000061000000600000005f",
        MEM_0D                  =>  x"0000006e0000006d0000006c0000006b0000006a000000690000006800000067",
        MEM_0E                  =>  x"000000760000007500000074000000730000007200000071000000700000006f",
        MEM_0F                  =>  x"0000007e0000007d0000007c0000007b0000007a000000790000007800000077",
        MEM_10                  =>  x"0000000600000005000000040000000300000002000000bc0000000100000000",
        MEM_11                  =>  x"0000000e0000000d0000000c0000000b0000000a000000090000000800000007",
        MEM_12                  =>  x"000000160000001500000014000000130000001200000011000000100000000f",
        MEM_13                  =>  x"0000001e0000001d0000001c0000001b0000001a000000190000001800000017",
        MEM_14                  =>  x"000000260000002500000024000000230000002200000021000000200000001f",
        MEM_15                  =>  x"0000002e0000002d0000002c0000002b0000002a000000290000002800000027",
        MEM_16                  =>  x"000000360000003500000034000000330000003200000031000000300000002f",
        MEM_17                  =>  x"0000003e0000003d0000003c0000003b0000003a000000390000003800000037",
        MEM_18                  =>  x"000000460000004500000044000000430000004200000041000000400000003f",
        MEM_19                  =>  x"0000004e0000004d0000004c0000004b0000004a000000490000004800000047",
        MEM_1A                  =>  x"000000560000005500000054000000530000005200000051000000500000004f",
        MEM_1B                  =>  x"0000005e0000005d0000005c0000005b0000005a000000590000005800000057",
        MEM_1C                  =>  x"000000660000006500000064000000630000006200000061000000600000005f",
        MEM_1D                  =>  x"0000006e0000006d0000006c0000006b0000006a000000690000006800000067",
        MEM_1E                  =>  x"000000760000007500000074000000730000007200000071000000700000006f",
        MEM_1F                  =>  x"0000007e0000007d0000007c0000007b0000007a000000790000007800000077",
        MEM_20                  =>  x"0000000600000005000000040000000300000002000000bc0000000100000000",
        MEM_21                  =>  x"0000000e0000000d0000000c0000000b0000000a000000090000000800000007",
        MEM_22                  =>  x"000000160000001500000014000000130000001200000011000000100000000f",
        MEM_23                  =>  x"0000001e0000001d0000001c0000001b0000001a000000190000001800000017",
        MEM_24                  =>  x"000000260000002500000024000000230000002200000021000000200000001f",
        MEM_25                  =>  x"0000002e0000002d0000002c0000002b0000002a000000290000002800000027",
        MEM_26                  =>  x"000000360000003500000034000000330000003200000031000000300000002f",
        MEM_27                  =>  x"0000003e0000003d0000003c0000003b0000003a000000390000003800000037",
        MEM_28                  =>  x"000000460000004500000044000000430000004200000041000000400000003f",
        MEM_29                  =>  x"0000004e0000004d0000004c0000004b0000004a000000490000004800000047",
        MEM_2A                  =>  x"000000560000005500000054000000530000005200000051000000500000004f",
        MEM_2B                  =>  x"0000005e0000005d0000005c0000005b0000005a000000590000005800000057",
        MEM_2C                  =>  x"000000660000006500000064000000630000006200000061000000600000005f",
        MEM_2D                  =>  x"0000006e0000006d0000006c0000006b0000006a000000690000006800000067",
        MEM_2E                  =>  x"000000760000007500000074000000730000007200000071000000700000006f",
        MEM_2F                  =>  x"0000007e0000007d0000007c0000007b0000007a000000790000007800000077",
        MEM_30                  =>  x"0000000600000005000000040000000300000002000000bc0000000100000000",
        MEM_31                  =>  x"0000000e0000000d0000000c0000000b0000000a000000090000000800000007",
        MEM_32                  =>  x"000000160000001500000014000000130000001200000011000000100000000f",
        MEM_33                  =>  x"0000001e0000001d0000001c0000001b0000001a000000190000001800000017",
        MEM_34                  =>  x"000000260000002500000024000000230000002200000021000000200000001f",
        MEM_35                  =>  x"0000002e0000002d0000002c0000002b0000002a000000290000002800000027",
        MEM_36                  =>  x"000000360000003500000034000000330000003200000031000000300000002f",
        MEM_37                  =>  x"0000003e0000003d0000003c0000003b0000003a000000390000003800000037",
        MEM_38                  =>  x"000000460000004500000044000000430000004200000041000000400000003f",
        MEM_39                  =>  x"0000004e0000004d0000004c0000004b0000004a000000490000004800000047",
        MEM_3A                  =>  x"000000560000005500000054000000530000005200000051000000500000004f",
        MEM_3B                  =>  x"0000005e0000005d0000005c0000005b0000005a000000590000005800000057",
        MEM_3C                  =>  x"000000660000006500000064000000630000006200000061000000600000005f",
        MEM_3D                  =>  x"0000006e0000006d0000006c0000006b0000006a000000690000006800000067",
        MEM_3E                  =>  x"000000760000007500000074000000730000007200000071000000700000006f",
        MEM_3F                  =>  x"0000007e0000007d0000007c0000007b0000007a000000790000007800000077",
        MEMP_00                  =>  x"0000000000000000000000000000000000000000000000000000000000000100",
        MEMP_01                  =>  x"0000000000000000000000000000000000000000000000000000000000000000",
        MEMP_02                  =>  x"0000000000000000000000000000000000000000000000000000000000000100",
        MEMP_03                  =>  x"0000000000000000000000000000000000000000000000000000000000000000",
        MEMP_04                  =>  x"0000000000000000000000000000000000000000000000000000000000000100",
        MEMP_05                  =>  x"0000000000000000000000000000000000000000000000000000000000000000",
        MEMP_06                  =>  x"0000000000000000000000000000000000000000000000000000000000000100",
        MEMP_07                  =>  x"0000000000000000000000000000000000000000000000000000000000000000"
    )
    port map
    (
        -- MGT Interface
        RX_DATA                         =>      tile0_rxdata0_i,
        RX_ENMCOMMA_ALIGN               =>      tile0_rxenmcommaalign0_i,
        RX_ENPCOMMA_ALIGN               =>      tile0_rxenpcommaalign0_i,
        RX_ENCHAN_SYNC                  =>      open,
        RX_CHANBOND_SEQ                 =>      tied_to_ground_i,
        -- Control Interface
        INC_IN                          =>      tile0_inc_in0_i,
        INC_OUT                         =>      tile0_inc_out0_i,
        PATTERN_MATCH_N                 =>      tile0_matchn0_i,
        RESET_ON_ERROR                  =>      tile0_frame_check0_reset_i,
        -- System Interface
        USER_CLK                        =>      tile0_txusrclk0_i,
        SYSTEM_RESET                    =>      tile0_rx_system_reset0_c,
        ERROR_COUNT                     =>      tile0_error_count0_i,
        TRACK_DATA                      =>      tile0_track_data0_i
    );
    
    tile0_frame_check1_reset_i              <= reset_on_data_error_i when (EXAMPLE_CONFIG_INDEPENDENT_LANES=0) else tile0_matchn1_i;

    -- tile0_frame_check0 is always connected to the lane with the start of char
    -- and this lane starts off the data checking on all the other lanes. The INC_IN port is tied off
    tile0_inc_in1_i                         <= '0';

    tile0_frame_check1 : FRAME_CHECK
    generic map
    (
        RX_DATA_WIDTH                   =>      8,
        USE_COMMA                       =>      1,
        WORDS_IN_BRAM                   =>      EXAMPLE_WORDS_IN_BRAM,
        CONFIG_INDEPENDENT_LANES        =>      1,
        START_OF_PACKET_CHAR            =>      x"bc",
        MEM_00                  =>  x"0000000600000005000000040000000300000002000000bc0000000100000000",
        MEM_01                  =>  x"0000000e0000000d0000000c0000000b0000000a000000090000000800000007",
        MEM_02                  =>  x"000000160000001500000014000000130000001200000011000000100000000f",
        MEM_03                  =>  x"0000001e0000001d0000001c0000001b0000001a000000190000001800000017",
        MEM_04                  =>  x"000000260000002500000024000000230000002200000021000000200000001f",
        MEM_05                  =>  x"0000002e0000002d0000002c0000002b0000002a000000290000002800000027",
        MEM_06                  =>  x"000000360000003500000034000000330000003200000031000000300000002f",
        MEM_07                  =>  x"0000003e0000003d0000003c0000003b0000003a000000390000003800000037",
        MEM_08                  =>  x"000000460000004500000044000000430000004200000041000000400000003f",
        MEM_09                  =>  x"0000004e0000004d0000004c0000004b0000004a000000490000004800000047",
        MEM_0A                  =>  x"000000560000005500000054000000530000005200000051000000500000004f",
        MEM_0B                  =>  x"0000005e0000005d0000005c0000005b0000005a000000590000005800000057",
        MEM_0C                  =>  x"000000660000006500000064000000630000006200000061000000600000005f",
        MEM_0D                  =>  x"0000006e0000006d0000006c0000006b0000006a000000690000006800000067",
        MEM_0E                  =>  x"000000760000007500000074000000730000007200000071000000700000006f",
        MEM_0F                  =>  x"0000007e0000007d0000007c0000007b0000007a000000790000007800000077",
        MEM_10                  =>  x"0000000600000005000000040000000300000002000000bc0000000100000000",
        MEM_11                  =>  x"0000000e0000000d0000000c0000000b0000000a000000090000000800000007",
        MEM_12                  =>  x"000000160000001500000014000000130000001200000011000000100000000f",
        MEM_13                  =>  x"0000001e0000001d0000001c0000001b0000001a000000190000001800000017",
        MEM_14                  =>  x"000000260000002500000024000000230000002200000021000000200000001f",
        MEM_15                  =>  x"0000002e0000002d0000002c0000002b0000002a000000290000002800000027",
        MEM_16                  =>  x"000000360000003500000034000000330000003200000031000000300000002f",
        MEM_17                  =>  x"0000003e0000003d0000003c0000003b0000003a000000390000003800000037",
        MEM_18                  =>  x"000000460000004500000044000000430000004200000041000000400000003f",
        MEM_19                  =>  x"0000004e0000004d0000004c0000004b0000004a000000490000004800000047",
        MEM_1A                  =>  x"000000560000005500000054000000530000005200000051000000500000004f",
        MEM_1B                  =>  x"0000005e0000005d0000005c0000005b0000005a000000590000005800000057",
        MEM_1C                  =>  x"000000660000006500000064000000630000006200000061000000600000005f",
        MEM_1D                  =>  x"0000006e0000006d0000006c0000006b0000006a000000690000006800000067",
        MEM_1E                  =>  x"000000760000007500000074000000730000007200000071000000700000006f",
        MEM_1F                  =>  x"0000007e0000007d0000007c0000007b0000007a000000790000007800000077",
        MEM_20                  =>  x"0000000600000005000000040000000300000002000000bc0000000100000000",
        MEM_21                  =>  x"0000000e0000000d0000000c0000000b0000000a000000090000000800000007",
        MEM_22                  =>  x"000000160000001500000014000000130000001200000011000000100000000f",
        MEM_23                  =>  x"0000001e0000001d0000001c0000001b0000001a000000190000001800000017",
        MEM_24                  =>  x"000000260000002500000024000000230000002200000021000000200000001f",
        MEM_25                  =>  x"0000002e0000002d0000002c0000002b0000002a000000290000002800000027",
        MEM_26                  =>  x"000000360000003500000034000000330000003200000031000000300000002f",
        MEM_27                  =>  x"0000003e0000003d0000003c0000003b0000003a000000390000003800000037",
        MEM_28                  =>  x"000000460000004500000044000000430000004200000041000000400000003f",
        MEM_29                  =>  x"0000004e0000004d0000004c0000004b0000004a000000490000004800000047",
        MEM_2A                  =>  x"000000560000005500000054000000530000005200000051000000500000004f",
        MEM_2B                  =>  x"0000005e0000005d0000005c0000005b0000005a000000590000005800000057",
        MEM_2C                  =>  x"000000660000006500000064000000630000006200000061000000600000005f",
        MEM_2D                  =>  x"0000006e0000006d0000006c0000006b0000006a000000690000006800000067",
        MEM_2E                  =>  x"000000760000007500000074000000730000007200000071000000700000006f",
        MEM_2F                  =>  x"0000007e0000007d0000007c0000007b0000007a000000790000007800000077",
        MEM_30                  =>  x"0000000600000005000000040000000300000002000000bc0000000100000000",
        MEM_31                  =>  x"0000000e0000000d0000000c0000000b0000000a000000090000000800000007",
        MEM_32                  =>  x"000000160000001500000014000000130000001200000011000000100000000f",
        MEM_33                  =>  x"0000001e0000001d0000001c0000001b0000001a000000190000001800000017",
        MEM_34                  =>  x"000000260000002500000024000000230000002200000021000000200000001f",
        MEM_35                  =>  x"0000002e0000002d0000002c0000002b0000002a000000290000002800000027",
        MEM_36                  =>  x"000000360000003500000034000000330000003200000031000000300000002f",
        MEM_37                  =>  x"0000003e0000003d0000003c0000003b0000003a000000390000003800000037",
        MEM_38                  =>  x"000000460000004500000044000000430000004200000041000000400000003f",
        MEM_39                  =>  x"0000004e0000004d0000004c0000004b0000004a000000490000004800000047",
        MEM_3A                  =>  x"000000560000005500000054000000530000005200000051000000500000004f",
        MEM_3B                  =>  x"0000005e0000005d0000005c0000005b0000005a000000590000005800000057",
        MEM_3C                  =>  x"000000660000006500000064000000630000006200000061000000600000005f",
        MEM_3D                  =>  x"0000006e0000006d0000006c0000006b0000006a000000690000006800000067",
        MEM_3E                  =>  x"000000760000007500000074000000730000007200000071000000700000006f",
        MEM_3F                  =>  x"0000007e0000007d0000007c0000007b0000007a000000790000007800000077",
        MEMP_00                  =>  x"0000000000000000000000000000000000000000000000000000000000000100",
        MEMP_01                  =>  x"0000000000000000000000000000000000000000000000000000000000000000",
        MEMP_02                  =>  x"0000000000000000000000000000000000000000000000000000000000000100",
        MEMP_03                  =>  x"0000000000000000000000000000000000000000000000000000000000000000",
        MEMP_04                  =>  x"0000000000000000000000000000000000000000000000000000000000000100",
        MEMP_05                  =>  x"0000000000000000000000000000000000000000000000000000000000000000",
        MEMP_06                  =>  x"0000000000000000000000000000000000000000000000000000000000000100",
        MEMP_07                  =>  x"0000000000000000000000000000000000000000000000000000000000000000"
    )
    port map
    (
        -- MGT Interface
        RX_DATA                         =>      tile0_rxdata1_i,
        RX_ENMCOMMA_ALIGN               =>      tile0_rxenmcommaalign1_i,
        RX_ENPCOMMA_ALIGN               =>      tile0_rxenpcommaalign1_i,
        RX_ENCHAN_SYNC                  =>      open,
        RX_CHANBOND_SEQ                 =>      tied_to_ground_i,
        -- Control Interface
        INC_IN                          =>      tile0_inc_in1_i,
        INC_OUT                         =>      tile0_inc_out1_i,
        PATTERN_MATCH_N                 =>      tile0_matchn1_i,
        RESET_ON_ERROR                  =>      tile0_frame_check1_reset_i,
        -- System Interface
        USER_CLK                        =>      tile0_txusrclk0_i,
        SYSTEM_RESET                    =>      tile0_rx_system_reset1_c,
        ERROR_COUNT                     =>      tile0_error_count1_i,
        TRACK_DATA                      =>      tile0_track_data1_i
    );
    

    TRACK_DATA_OUT                          <= track_data_out_i;

    track_data_out_i                        <= 
                                tile0_track_data0_i  and
                                tile0_track_data1_i ;


    reset_on_data_error_i                   <= '0';



    ----------------------------- Chipscope Connections -----------------------
    -- When the example design is run in hardware, it uses chipscope to allow the
    -- example design and GTP wrapper to be controlled and monitored. The 
    -- EXAMPLE_USE_CHIPSCOPE parameter allows chipscope to be removed for simulation.
    
chipscope : if EXAMPLE_USE_CHIPSCOPE = 1 generate


    -- Shared VIO for all tiles
    shared_vio_i : shared_vio
    port map
    (
        control                         =>      shared_vio_control_i,
        async_in                        =>      shared_vio_in_i,
        async_out                       =>      shared_vio_out_i
    );

    
    -- ICON for all VIOs 
    i_icon : icon
    port map
    (
        control0                        =>      shared_vio_control_i,
        control1                        =>      tile0_data_vio_control_i,
        control2                        =>      tile0_gtp0_ila_control_i,
        control3                        =>      tile0_gtp1_ila_control_i,
        control4                        =>      null_vio_4_i,
        control5                        =>      null_vio_5_i,
        control6                        =>      null_vio_6_i,
        control7                        =>      null_vio_7_i,
        control8                        =>      null_vio_8_i,
        control9                        =>      null_vio_9_i,
        control10                       =>      null_vio_10_i,
        control11                       =>      null_vio_11_i,
        control12                       =>      null_vio_12_i
    );

    -- TILE0 DATA VIO 
    tile0_data_vio_i : data_vio
    port map
    (
        control                         =>      tile0_data_vio_control_i,
        async_in                        =>      tile0_data_vio_in_i,
        async_out                       =>      tile0_data_vio_out_i    
    );
    
    -- TILE0 GTP0 RX ILA 
    tile0_gtp0_i : ila
    port map
    (
        control                         =>      tile0_gtp0_ila_control_i,
        clk                             =>      tile0_txusrclk0_i,
        trig0                           =>      tile0_ila_in0_i
    );
    -- TILE0 GTP1 RX ILA 
    tile0_gtp1_i : ila
    port map
    (
        control                         =>      tile0_gtp1_ila_control_i,
        clk                             =>      tile0_txusrclk0_i,
        trig0                           =>      tile0_ila_in1_i
    );
    


    i_null_vio_4 : null_vio
    port map
    (
        control                         =>      null_vio_4_i
    );
    
    i_null_vio_5 : null_vio
    port map
    (
        control                         =>      null_vio_5_i
    );
    
    i_null_vio_6 : null_vio
    port map
    (
        control                         =>      null_vio_6_i
    );
    
    i_null_vio_7 : null_vio
    port map
    (
        control                         =>      null_vio_7_i
    );
    
    i_null_vio_8 : null_vio
    port map
    (
        control                         =>      null_vio_8_i
    );
    
    i_null_vio_9 : null_vio
    port map
    (
        control                         =>      null_vio_9_i
    );
    
    i_null_vio_10 : null_vio
    port map
    (
        control                         =>      null_vio_10_i
    );
    
    i_null_vio_11 : null_vio
    port map
    (
        control                         =>      null_vio_11_i
    );
    
    i_null_vio_12 : null_vio
    port map
    (
        control                         =>      null_vio_12_i
    );
    


    -- Connect resets for frame generators
    tile0_tx_system_reset0_c                <= not tile0_tx_resetdone0_r2 or user_tx_reset_i;
    tile0_tx_system_reset1_c                <= not tile0_tx_resetdone1_r2 or user_tx_reset_i;
    tile0_rx_system_reset0_c                <= not tile0_rx_resetdone0_r2 or user_rx_reset_i;
    tile0_rx_system_reset1_c                <= not tile0_rx_resetdone1_r2 or user_rx_reset_i;


    tile0_gtpreset0_i                       <= gtpreset0_i;
    tile0_gtpreset1_i                       <= gtpreset0_i;   


    -- Shared VIO Outputs
    gtpreset0_i                             <= shared_vio_out_i(31);
    user_tx_reset_i                         <= shared_vio_out_i(30);
    user_rx_reset_i                         <= shared_vio_out_i(29);

    -- Shared VIO Inputs
    shared_vio_in_i(31)                     <= tile0_plllkdet0_i;
    shared_vio_in_i(30 downto 0)            <= tied_to_ground_vec_i(30 downto 0);

    -- Chipscope VIO input connections on Tile 0
    tile0_data_vio_in_i(139)                <= tile0_resetdone0_i;
    tile0_data_vio_in_i(138)                <= tile0_resetdone1_i;
    tile0_data_vio_in_i(137 downto 136)     <= tile0_txbufstatus0_i;
    tile0_data_vio_in_i(135 downto 134)     <= tile0_txbufstatus1_i;
    tile0_data_vio_in_i(133 downto 0)       <= tied_to_ground_vec_i(133 downto 0);

    -- Chipscope VIO ouptut connections on Tile 0
    tile0_loopback0_i                       <= tile0_data_vio_out_i(139 downto 137);
    tile0_loopback1_i                       <= tile0_data_vio_out_i(136 downto 134);
    tile0_rxpowerdown0_i                    <= tile0_data_vio_out_i(133 downto 132);
    tile0_rxpowerdown1_i                    <= tile0_data_vio_out_i(131 downto 130);
    tile0_txpowerdown0_i                    <= tile0_data_vio_out_i(129 downto 128);
    tile0_txpowerdown1_i                    <= tile0_data_vio_out_i(127 downto 126);
    tile0_rxbufreset0_i                     <= tile0_data_vio_out_i(125);
    tile0_rxbufreset1_i                     <= tile0_data_vio_out_i(124);
    tile0_txchardispmode0_i                 <= tile0_data_vio_out_i(123);
    tile0_txchardispmode1_i                 <= tile0_data_vio_out_i(122);
    tile0_txchardispval0_i                  <= tile0_data_vio_out_i(121);
    tile0_txchardispval1_i                  <= tile0_data_vio_out_i(120);

    -- Chipscope ILA connections for GTP0 on Tile 0
    tile0_ila_in0_i(84)                     <= tile0_rxchariscomma0_i;
    tile0_ila_in0_i(83)                     <= tile0_rxcharisk0_i;
    tile0_ila_in0_i(82)                     <= tile0_rxdisperr0_i;
    tile0_ila_in0_i(81)                     <= tile0_rxnotintable0_i;
    tile0_ila_in0_i(80)                     <= tile0_rxrundisp0_i;
    tile0_ila_in0_i(79 downto 77)           <= tile0_rxclkcorcnt0_i;
    tile0_ila_in0_i(76 downto 69)           <= tile0_rxdata0_i;
    tile0_ila_in0_i(68 downto 66)           <= tile0_rxbufstatus0_i;
    tile0_ila_in0_i(65 downto 58)           <= tile0_error_count0_i;
    tile0_ila_in0_i(57 downto 0)            <= tied_to_ground_vec_i(57 downto 0);

    -- Chipscope ILA connections for GTP1 on Tile 0
    tile0_ila_in1_i(84)                     <= tile0_rxchariscomma1_i;
    tile0_ila_in1_i(83)                     <= tile0_rxcharisk1_i;
    tile0_ila_in1_i(82)                     <= tile0_rxdisperr1_i;
    tile0_ila_in1_i(81)                     <= tile0_rxnotintable1_i;
    tile0_ila_in1_i(80)                     <= tile0_rxrundisp1_i;
    tile0_ila_in1_i(79 downto 77)           <= tile0_rxclkcorcnt1_i;
    tile0_ila_in1_i(76 downto 69)           <= tile0_rxdata1_i;
    tile0_ila_in1_i(68 downto 66)           <= tile0_rxbufstatus1_i;
    tile0_ila_in1_i(65 downto 58)           <= tile0_error_count1_i;
    tile0_ila_in1_i(57 downto 0)            <= tied_to_ground_vec_i(57 downto 0);


   
end generate chipscope;


no_chipscope : if EXAMPLE_USE_CHIPSCOPE = 0 generate

    -- If Chipscope is not being used, drive GTP reset signal
    -- from the top level ports
    tile0_gtpreset0_i                       <= GTP0_RESET_IN;
    tile0_gtpreset1_i                       <= GTP1_RESET_IN;

    -- assign resets for frame_gen and frame_check modules
    tile0_tx_system_reset0_c                <= not tile0_tx_resetdone0_r2;
    tile0_tx_system_reset1_c                <= not tile0_tx_resetdone1_r2;
    tile0_rx_system_reset0_c                <= not tile0_rx_resetdone0_r2;
    tile0_rx_system_reset1_c                <= not tile0_rx_resetdone1_r2;

    gtpreset0_i                             <= tied_to_ground_i;
    user_tx_reset_i                         <= tied_to_ground_i;
    user_rx_reset_i                         <= tied_to_ground_i;
    tile0_loopback0_i                       <= tied_to_ground_vec_i(2 downto 0);
    tile0_loopback1_i                       <= tied_to_ground_vec_i(2 downto 0);
    tile0_rxpowerdown0_i                    <= tied_to_ground_vec_i(1 downto 0);
    tile0_rxpowerdown1_i                    <= tied_to_ground_vec_i(1 downto 0);
    tile0_txpowerdown0_i                    <= tied_to_ground_vec_i(1 downto 0);
    tile0_txpowerdown1_i                    <= tied_to_ground_vec_i(1 downto 0);
    tile0_rxbufreset0_i                     <= tied_to_ground_i;
    tile0_rxbufreset1_i                     <= tied_to_ground_i;
    tile0_txchardispmode0_i                 <= tied_to_ground_i;
    tile0_txchardispmode1_i                 <= tied_to_ground_i;
    tile0_txchardispval0_i                  <= tied_to_ground_i;
    tile0_txchardispval1_i                  <= tied_to_ground_i;



end generate no_chipscope;


end RTL;

